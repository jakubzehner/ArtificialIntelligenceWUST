module main

import reversi
import ai

fn main() {
	// reversi.test()
	ai.test()
}
