module main

import reversi

fn main() {
	reversi.test()
}
