module reversi

pub struct Move {
pub:
	x int
	y int
}
