module reversi

pub enum Result {
	white_winner
	black_winner
	draw
}
